module Datapath(
ALUop,
MemtoReg,
MemRead,
MemWrite,
IorD,
RegWrite,
ALuSrc,
CLOCK_50);

input [3:0] ALUop;


endmodule