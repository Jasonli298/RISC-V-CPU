module seg7(
input [3:0] in,
input en,
output [6:0] HEX);



endmodule
